module up_counter(
    input  wire clk,
    input  wire rst,      // synchronous reset
    output reg  [2:0] q
);

always @(posedge clk) begin
    if (rst)
        q <= 3'b000;
    else
        q <= q + 1'b1;
end

endmodule